// Syndrome → Coset Leader LUT (hardcoded to match python_simulation COSET_LEADERS)
module coset_leader_lut (
    input  wire [5:0] syndrome,      // 6-bit key (tuple order: row0..row5)
    output reg  [12:0] leader        // 13-bit coset leader (v bits)
);
    // Address packs syndrome bits in tuple order: {row0,row1,row2,row3,row4,row5}
    wire [5:0] addr = {syndrome[0], syndrome[1], syndrome[2], syndrome[3], syndrome[4], syndrome[5]};

    // Mapping: python index i (0..12) → Verilog bit (12-i)
    // So a python vector with 1 at index 0 becomes 13'b1000000000000, index 12 → 13'b0000000000001
    always @* begin
        case (addr)
            6'b000000: leader = 13'b0000000000000; // (0,0,0,0,0,0)
            6'b100000: leader = 13'b1000000000000; // (1,0,0,0,0,0)
            6'b010000: leader = 13'b0100000000000; // (0,1,0,0,0,0)
            6'b110000: leader = 13'b1100000000000; // (1,1,0,0,0,0)
            6'b001000: leader = 13'b0010000000000; // (0,0,1,0,0,0)
            6'b101000: leader = 13'b1010000000000; // (1,0,1,0,0,0)
            6'b011000: leader = 13'b0110000000000; // (0,1,1,0,0,0)
            6'b111000: leader = 13'b0000001000010; // (1,1,1,0,0,0)
            6'b000100: leader = 13'b0001000000000; // (0,0,0,1,0,0)
            6'b100100: leader = 13'b1001000000000; // (1,0,0,1,0,0)
            6'b010100: leader = 13'b0101000000000; // (0,1,0,1,0,0)
            6'b110100: leader = 13'b0000000001100; // (1,1,0,1,0,0)
            6'b001100: leader = 13'b0011000000000; // (0,0,1,1,0,0)
            6'b101100: leader = 13'b0000000001001; // (1,0,1,1,0,0)
            6'b011100: leader = 13'b0000100001000; // (0,1,1,1,0,0)
            6'b111100: leader = 13'b0000001100000; // (1,1,1,1,0,0)
            6'b000010: leader = 13'b0000100000000; // (0,0,0,0,1,0)
            6'b100010: leader = 13'b1000100000000; // (1,0,0,0,1,0)
            6'b010010: leader = 13'b0100100000000; // (0,1,0,0,1,0)
            6'b110010: leader = 13'b0000010100000; // (1,1,0,0,1,0)
            6'b001010: leader = 13'b0010100000000; // (0,0,1,0,1,0)
            6'b101010: leader = 13'b0000000001000; // (1,0,1,0,1,0) matches Python index 9
            6'b011010: leader = 13'b0000010100000; // (0,1,1,0,1,0)
            6'b111010: leader = 13'b0100000100000; // (1,1,1,0,1,0)
            6'b000110: leader = 13'b0001100000000; // (0,0,0,1,1,0)
            6'b100110: leader = 13'b0000001100000; // (1,0,0,1,1,0)
            6'b010110: leader = 13'b0010000100000; // (0,1,0,1,1,0)
            6'b110110: leader = 13'b0000001000010; // (1,1,0,1,1,0)
            6'b001110: leader = 13'b0000110000000; // (0,0,1,1,1,0)
            6'b101110: leader = 13'b0000100001000; // (1,0,1,1,1,0)
            6'b011110: leader = 13'b0000000001000; // (0,1,1,1,1,0)
            6'b111110: leader = 13'b1000000001000; // (1,1,1,1,1,0)
            6'b000001: leader = 13'b0000010000000; // (0,0,0,0,0,1)
            6'b100001: leader = 13'b1000010000000; // (1,0,0,0,0,1)
            6'b010001: leader = 13'b0100010000000; // (0,1,0,0,0,1)
            6'b110001: leader = 13'b0000100100000; // (1,1,0,0,0,1)
            6'b001001: leader = 13'b0010010000000; // (0,0,1,0,0,1)
            6'b101001: leader = 13'b0100000000010; // (1,0,1,0,0,1)
            6'b011001: leader = 13'b0000010101000; // (0,1,1,0,0,1)
            6'b111001: leader = 13'b0000000000010; // (1,1,1,0,0,1)
            6'b000101: leader = 13'b0001010000000; // (0,0,0,1,0,1)
            6'b100101: leader = 13'b0001001001000; // (1,0,0,1,0,1)
            6'b010101: leader = 13'b0000000010000; // (0,1,0,1,0,1)
            6'b110101: leader = 13'b1000000100000; // (1,1,0,1,0,1)
            6'b001101: leader = 13'b0001011000000; // (0,0,1,1,0,1)
            6'b101101: leader = 13'b0000100100000; // (1,0,1,1,0,1)
            6'b011101: leader = 13'b0000000100000; // (0,1,1,1,0,1)
            6'b111101: leader = 13'b1000001000000; // (1,1,1,1,0,1)
            6'b000011: leader = 13'b0000110000000; // (0,0,0,0,1,1)
            6'b100011: leader = 13'b0100010001000; // (1,0,0,0,1,1)
            6'b010011: leader = 13'b1000010001000; // (0,1,0,0,1,1)
            6'b110011: leader = 13'b0000010000000; // (1,1,0,0,1,1)
            6'b001011: leader = 13'b0001010000000; // (0,0,1,0,1,1)
            6'b101011: leader = 13'b0000100010000; // (1,0,1,0,1,1)
            6'b011011: leader = 13'b0000000000001; // (0,1,1,0,1,1)
            6'b111011: leader = 13'b0010001000000; // (1,1,1,0,1,1)
            6'b000111: leader = 13'b0010010000000; // (0,0,0,1,1,1)
            6'b100111: leader = 13'b0000000001100; // (1,0,0,1,1,1)
            6'b010111: leader = 13'b0000100010000; // (0,1,0,1,1,1)
            6'b110111: leader = 13'b0001000100000; // (1,1,0,1,1,1)
            6'b001111: leader = 13'b0000001000000; // (0,0,1,1,1,1)
            6'b101111: leader = 13'b1000001000000; // (1,0,1,1,1,1)
            6'b011111: leader = 13'b0100001000000; // (0,1,1,1,1,1)
            6'b111111: leader = 13'b0000001100000; // (1,1,1,1,1,1)
            default:   leader = 13'b0000000000000;
        endcase
    end
endmodule


