`timescale 1 ns / 1 ps
module sakura_g_main_ring_osc_tb;

	parameter symbol_time = 17361.1;

	reg clk;
	reg rst_n;
	reg rx;
	wire tx;
	wire M_HEADER;	
	wire M_LED_0;	

	
	sakura_g_main_ring_osc // PUT YOUR TOP LEVEL (WITH/WITHOUT PLL)
	dut (
		.M_CLK_OSC    (clk),
		.M_RESET_B    (rst_n),
		.FTDI_BDBUS_0 (rx),
		.FTDI_BDBUS_1 (tx),
		.M_HEADER     (M_HEADER),
		.M_LED_0 	  (M_LED_0),
		.M_LED_1      ()
	);

	task send_uart_byte; // TASK THAT RECEIVES A BYTE AND SENDS IT SERIALLY VIA UART
		input [7:0] in_byte;
	begin 
		//$display("sending byte %0h", in_byte);
		repeat (4) @(posedge clk);
		#(symbol_time) rx = 1'b0; // start bit
		#(symbol_time) rx = in_byte[0];
		#(symbol_time) rx = in_byte[1];
		#(symbol_time) rx = in_byte[2];
		#(symbol_time) rx = in_byte[3];
		#(symbol_time) rx = in_byte[4];
		#(symbol_time) rx = in_byte[5];
		#(symbol_time) rx = in_byte[6];
		#(symbol_time) rx = in_byte[7];
		#(symbol_time) rx = 1'b1; // stop bit
		repeat (4) @(posedge clk);
		repeat (40) @(posedge clk);

	end
	endtask

	always #(20.8333/2) clk = ~clk; //48MHZ clock (IF USING PLL)
	//always #(250/2) clk = ~clk;     //4MHZ clock (IF NOT USING PLL)

	initial begin
		clk = 0;
		rst_n = 0;
		rx = 1;
		repeat (4) @(posedge clk);

		rst_n = 1;
	
		send_uart_byte(8'h00);
		send_uart_byte(8'h00);
		
		send_uart_byte(8'hFF);
		send_uart_byte(8'hFF);
		
		send_uart_byte(8'h00);
		send_uart_byte(8'h00);
	
		repeat (100000) @(posedge clk);

		$finish;


	end
endmodule
